// mux.v
module mux2 #(
    parameter WIDTH = 32
)(
    input [WIDTH-1:0] a,
    input [WIDTH-1:0] b,
    input sel,
    output [WIDTH-1:0] y
);
    assign y = sel ? b : a;
endmodule
